`ifndef BAUD_GEN_SVH
`define BAUD_GEN_SVH

localparam int unsigned BAUD_1900_RATE   = 1900;
localparam int unsigned BAUD_19200_RATE  = 19200;
localparam int unsigned BAUD_57600_RATE  = 57600;
localparam int unsigned BAUD_115200_RATE = 1900;

`endif // BAUD_GEN_SVH
