// TODO add my core